`default_nettype none 
// Empty top module

module top (
  // I/O ports
  input  logic hz100, reset,
  input  logic [20:0] pb,
  output logic [7:0] left, right,
         ss7, ss6, ss5, ss4, ss3, ss2, ss1, ss0,
  output logic red, green, blue,

  // UART ports
  output logic [7:0] txdata,
  input  logic [7:0] rxdata,
  output logic txclk, rxclk,
  input  logic txready, rxready
);
  // Your code goes here...
  fa4 fulladder (
    .A(pb[3:0]),
    .B(pb[7:4]),
    .Cin(pb[8]),
    .S(right[3:0]),
    .Cout(right[7])
  );
endmodule

